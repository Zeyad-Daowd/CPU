library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
use std.textio.all;
use ieee.std_logic_textio.all;

entity Instruction_Memory is
    port (
        clk: in std_logic; -- Clock 
        -- for reading the instructions
        pc: in std_logic_vector(15 downto 0); -- read address [PC]
        instruction: out std_logic_vector(15 downto 0); -- 16-bit instruction 
        -- for writing the instructions
        write_enable: in std_logic;  -- Write enable signal
        write_address: in std_logic_vector(15 downto 0); -- 16-bit write address, like pc
        write_data: in std_logic_vector(15 downto 0) -- 16-bit instruction to be written
    );
end Instruction_Memory;

architecture Behavioral of Instruction_Memory is
    -- memory array
    type memory_array is array (0 to 4095) of std_logic_vector(15 downto 0);
    
    
    signal memory: memory_array := (
        0 => "0000011100000000",
        1 => "0000010000000000",
        2 => "0000011000000000",
        3 => "0000000000000000",
        4 => "0000000000000000",
        5 => "0000000000000000",
        6 => "0000100000000000",
        7 => "0000000000000000",
        8 => "0000101000000000",
        9 => "0000000000000000",
        10 => "0000000000000000",
        11 => "0000000000000000",
        12 => "0000000000000000",
        13 => "0000000000000000",
        14 => "0000000000000000",
        15 => "0000000000000000",
        16 => "0000000000000000",
        17 => "0000000000000000",
        18 => "0000000000000000",
        19 => "0000000000000000",
        20 => "0000000000000000",
        21 => "0000000000000000",
        22 => "0000000000000000",
        23 => "0000000000000000",
        24 => "0000000000000000",
        25 => "0000000000000000",
        26 => "0000000000000000",
        27 => "0000000000000000",
        28 => "0000000000000000",
        29 => "0000000000000000",
        30 => "0000000000000000",
        31 => "0000000000000000",
        32 => "0000000000000000",
        33 => "0000000000000000",
        34 => "0000000000000000",
        35 => "0000000000000000",
        36 => "0000000000000000",
        37 => "0000000000000000",
        38 => "0000000000000000",
        39 => "0000000000000000",
        40 => "0000000000000000",
        41 => "0000000000000000",
        42 => "0000000000000000",
        43 => "0000000000000000",
        44 => "0000000000000000",
        45 => "0000000000000000",
        46 => "0000000000000000",
        47 => "0000000000000000",
        48 => "0101110100110100",
        49 => "1111000000000000",
        50 => "1100000001000000",
        51 => "0010011111100000",
        52 => "0000000000000000",
        53 => "0000000000000000",
        54 => "0000000000000000",
        55 => "0000000000000000",
        56 => "0000000000000000",
        57 => "0000000000000000",
        58 => "0000000000000000",
        59 => "0000000000000000",
        60 => "0000000000000000",
        61 => "0000000000000000",
        62 => "0000000000000000",
        63 => "0000000000000000",
        64 => "0000000000000000",
        65 => "0000000000000000",
        66 => "0000000000000000",
        67 => "0000000000000000",
        68 => "0000000000000000",
        69 => "0000000000000000",
        70 => "0000000000000000",
        71 => "0000000000000000",
        72 => "0000000000000000",
        73 => "0000000000000000",
        74 => "0000000000000000",
        75 => "0000000000000000",
        76 => "0000000000000000",
        77 => "0000000000000000",
        78 => "0000000000000000",
        79 => "0000000000000000",
        80 => "1100000001100000",
        81 => "0001110110100000",
        82 => "0010010110100000",
        83 => "0011011000000000",
        84 => "1100000011000000",
        85 => "0010000100100000",
        86 => "0000000000000000",
        87 => "0000000000000000",
        88 => "0000000000000000",
        89 => "0000000000000000",
        90 => "0000000000000000",
        91 => "0000000000000000",
        92 => "0000000000000000",
        93 => "0000000000000000",
        94 => "0000000000000000",
        95 => "0000000000000000",
        96 => "0000000000000000",
        97 => "0000000000000000",
        98 => "0000000000000000",
        99 => "0000000000000000",
        100 => "0000000000000000",
        101 => "0000000000000000",
        102 => "0000000000000000",
        103 => "0000000000000000",
        104 => "0000000000000000",
        105 => "0000000000000000",
        106 => "0000000000000000",
        107 => "0000000000000000",
        108 => "0000000000000000",
        109 => "0000000000000000",
        110 => "0000000000000000",
        111 => "0000000000000000",
        112 => "0000000000000000",
        113 => "0000000000000000",
        114 => "0000000000000000",
        115 => "0000000000000000",
        116 => "0000000000000000",
        117 => "0000000000000000",
        118 => "0000000000000000",
        119 => "0000000000000000",
        120 => "0000000000000000",
        121 => "0000000000000000",
        122 => "0000000000000000",
        123 => "0000000000000000",
        124 => "0000000000000000",
        125 => "0000000000000000",
        126 => "0000000000000000",
        127 => "0000000000000000",
        128 => "0000000000000000",
        129 => "0000000000000000",
        130 => "0000000000000000",
        131 => "0000000000000000",
        132 => "0000000000000000",
        133 => "0000000000000000",
        134 => "0000000000000000",
        135 => "0000000000000000",
        136 => "0000000000000000",
        137 => "0000000000000000",
        138 => "0000000000000000",
        139 => "0000000000000000",
        140 => "0000000000000000",
        141 => "0000000000000000",
        142 => "0000000000000000",
        143 => "0000000000000000",
        144 => "0000000000000000",
        145 => "0000000000000000",
        146 => "0000000000000000",
        147 => "0000000000000000",
        148 => "0000000000000000",
        149 => "0000000000000000",
        150 => "0000000000000000",
        151 => "0000000000000000",
        152 => "0000000000000000",
        153 => "0000000000000000",
        154 => "0000000000000000",
        155 => "0000000000000000",
        156 => "0000000000000000",
        157 => "0000000000000000",
        158 => "0000000000000000",
        159 => "0000000000000000",
        160 => "0000000000000000",
        161 => "0000000000000000",
        162 => "0000000000000000",
        163 => "0000000000000000",
        164 => "0000000000000000",
        165 => "0000000000000000",
        166 => "0000000000000000",
        167 => "0000000000000000",
        168 => "0000000000000000",
        169 => "0000000000000000",
        170 => "0000000000000000",
        171 => "0000000000000000",
        172 => "0000000000000000",
        173 => "0000000000000000",
        174 => "0000000000000000",
        175 => "0000000000000000",
        176 => "0000000000000000",
        177 => "0000000000000000",
        178 => "0000000000000000",
        179 => "0000000000000000",
        180 => "0000000000000000",
        181 => "0000000000000000",
        182 => "0000000000000000",
        183 => "0000000000000000",
        184 => "0000000000000000",
        185 => "0000000000000000",
        186 => "0000000000000000",
        187 => "0000000000000000",
        188 => "0000000000000000",
        189 => "0000000000000000",
        190 => "0000000000000000",
        191 => "0000000000000000",
        192 => "0000000000000000",
        193 => "0000000000000000",
        194 => "0000000000000000",
        195 => "0000000000000000",
        196 => "0000000000000000",
        197 => "0000000000000000",
        198 => "0000000000000000",
        199 => "0000000000000000",
        200 => "0000000000000000",
        201 => "0000000000000000",
        202 => "0000000000000000",
        203 => "0000000000000000",
        204 => "0000000000000000",
        205 => "0000000000000000",
        206 => "0000000000000000",
        207 => "0000000000000000",
        208 => "0000000000000000",
        209 => "0000000000000000",
        210 => "0000000000000000",
        211 => "0000000000000000",
        212 => "0000000000000000",
        213 => "0000000000000000",
        214 => "0000000000000000",
        215 => "0000000000000000",
        216 => "0000000000000000",
        217 => "0000000000000000",
        218 => "0000000000000000",
        219 => "0000000000000000",
        220 => "0000000000000000",
        221 => "0000000000000000",
        222 => "0000000000000000",
        223 => "0000000000000000",
        224 => "0000000000000000",
        225 => "0000000000000000",
        226 => "0000000000000000",
        227 => "0000000000000000",
        228 => "0000000000000000",
        229 => "0000000000000000",
        230 => "0000000000000000",
        231 => "0000000000000000",
        232 => "0000000000000000",
        233 => "0000000000000000",
        234 => "0000000000000000",
        235 => "0000000000000000",
        236 => "0000000000000000",
        237 => "0000000000000000",
        238 => "0000000000000000",
        239 => "0000000000000000",
        240 => "0000000000000000",
        241 => "0000000000000000",
        242 => "0000000000000000",
        243 => "0000000000000000",
        244 => "0000000000000000",
        245 => "0000000000000000",
        246 => "0000000000000000",
        247 => "0000000000000000",
        248 => "0000000000000000",
        249 => "0000000000000000",
        250 => "0000000000000000",
        251 => "0000000000000000",
        252 => "0000000000000000",
        253 => "0000000000000000",
        254 => "0000000000000000",
        255 => "0000000000000000",
        256 => "0000000000000000",
        257 => "0000000000000000",
        258 => "0000000000000000",
        259 => "0000000000000000",
        260 => "0000000000000000",
        261 => "0000000000000000",
        262 => "0000000000000000",
        263 => "0000000000000000",
        264 => "0000000000000000",
        265 => "0000000000000000",
        266 => "0000000000000000",
        267 => "0000000000000000",
        268 => "0000000000000000",
        269 => "0000000000000000",
        270 => "0000000000000000",
        271 => "0000000000000000",
        272 => "0000000000000000",
        273 => "0000000000000000",
        274 => "0000000000000000",
        275 => "0000000000000000",
        276 => "0000000000000000",
        277 => "0000000000000000",
        278 => "0000000000000000",
        279 => "0000000000000000",
        280 => "0000000000000000",
        281 => "0000000000000000",
        282 => "0000000000000000",
        283 => "0000000000000000",
        284 => "0000000000000000",
        285 => "0000000000000000",
        286 => "0000000000000000",
        287 => "0000000000000000",
        288 => "0000000000000000",
        289 => "0000000000000000",
        290 => "0000000000000000",
        291 => "0000000000000000",
        292 => "0000000000000000",
        293 => "0000000000000000",
        294 => "0000000000000000",
        295 => "0000000000000000",
        296 => "0000000000000000",
        297 => "0000000000000000",
        298 => "0000000000000000",
        299 => "0000000000000000",
        300 => "0000000000000000",
        301 => "0000000000000000",
        302 => "0000000000000000",
        303 => "0000000000000000",
        304 => "0000000000000000",
        305 => "0000000000000000",
        306 => "0000000000000000",
        307 => "0000000000000000",
        308 => "0000000000000000",
        309 => "0000000000000000",
        310 => "0000000000000000",
        311 => "0000000000000000",
        312 => "0000000000000000",
        313 => "0000000000000000",
        314 => "0000000000000000",
        315 => "0000000000000000",
        316 => "0000000000000000",
        317 => "0000000000000000",
        318 => "0000000000000000",
        319 => "0000000000000000",
        320 => "0000000000000000",
        321 => "0000000000000000",
        322 => "0000000000000000",
        323 => "0000000000000000",
        324 => "0000000000000000",
        325 => "0000000000000000",
        326 => "0000000000000000",
        327 => "0000000000000000",
        328 => "0000000000000000",
        329 => "0000000000000000",
        330 => "0000000000000000",
        331 => "0000000000000000",
        332 => "0000000000000000",
        333 => "0000000000000000",
        334 => "0000000000000000",
        335 => "0000000000000000",
        336 => "0000000000000000",
        337 => "0000000000000000",
        338 => "0000000000000000",
        339 => "0000000000000000",
        340 => "0000000000000000",
        341 => "0000000000000000",
        342 => "0000000000000000",
        343 => "0000000000000000",
        344 => "0000000000000000",
        345 => "0000000000000000",
        346 => "0000000000000000",
        347 => "0000000000000000",
        348 => "0000000000000000",
        349 => "0000000000000000",
        350 => "0000000000000000",
        351 => "0000000000000000",
        352 => "0000000000000000",
        353 => "0000000000000000",
        354 => "0000000000000000",
        355 => "0000000000000000",
        356 => "0000000000000000",
        357 => "0000000000000000",
        358 => "0000000000000000",
        359 => "0000000000000000",
        360 => "0000000000000000",
        361 => "0000000000000000",
        362 => "0000000000000000",
        363 => "0000000000000000",
        364 => "0000000000000000",
        365 => "0000000000000000",
        366 => "0000000000000000",
        367 => "0000000000000000",
        368 => "0000000000000000",
        369 => "0000000000000000",
        370 => "0000000000000000",
        371 => "0000000000000000",
        372 => "0000000000000000",
        373 => "0000000000000000",
        374 => "0000000000000000",
        375 => "0000000000000000",
        376 => "0000000000000000",
        377 => "0000000000000000",
        378 => "0000000000000000",
        379 => "0000000000000000",
        380 => "0000000000000000",
        381 => "0000000000000000",
        382 => "0000000000000000",
        383 => "0000000000000000",
        384 => "0000000000000000",
        385 => "0000000000000000",
        386 => "0000000000000000",
        387 => "0000000000000000",
        388 => "0000000000000000",
        389 => "0000000000000000",
        390 => "0000000000000000",
        391 => "0000000000000000",
        392 => "0000000000000000",
        393 => "0000000000000000",
        394 => "0000000000000000",
        395 => "0000000000000000",
        396 => "0000000000000000",
        397 => "0000000000000000",
        398 => "0000000000000000",
        399 => "0000000000000000",
        400 => "0000000000000000",
        401 => "0000000000000000",
        402 => "0000000000000000",
        403 => "0000000000000000",
        404 => "0000000000000000",
        405 => "0000000000000000",
        406 => "0000000000000000",
        407 => "0000000000000000",
        408 => "0000000000000000",
        409 => "0000000000000000",
        410 => "0000000000000000",
        411 => "0000000000000000",
        412 => "0000000000000000",
        413 => "0000000000000000",
        414 => "0000000000000000",
        415 => "0000000000000000",
        416 => "0000000000000000",
        417 => "0000000000000000",
        418 => "0000000000000000",
        419 => "0000000000000000",
        420 => "0000000000000000",
        421 => "0000000000000000",
        422 => "0000000000000000",
        423 => "0000000000000000",
        424 => "0000000000000000",
        425 => "0000000000000000",
        426 => "0000000000000000",
        427 => "0000000000000000",
        428 => "0000000000000000",
        429 => "0000000000000000",
        430 => "0000000000000000",
        431 => "0000000000000000",
        432 => "0000000000000000",
        433 => "0000000000000000",
        434 => "0000000000000000",
        435 => "0000000000000000",
        436 => "0000000000000000",
        437 => "0000000000000000",
        438 => "0000000000000000",
        439 => "0000000000000000",
        440 => "0000000000000000",
        441 => "0000000000000000",
        442 => "0000000000000000",
        443 => "0000000000000000",
        444 => "0000000000000000",
        445 => "0000000000000000",
        446 => "0000000000000000",
        447 => "0000000000000000",
        448 => "0000000000000000",
        449 => "0000000000000000",
        450 => "0000000000000000",
        451 => "0000000000000000",
        452 => "0000000000000000",
        453 => "0000000000000000",
        454 => "0000000000000000",
        455 => "0000000000000000",
        456 => "0000000000000000",
        457 => "0000000000000000",
        458 => "0000000000000000",
        459 => "0000000000000000",
        460 => "0000000000000000",
        461 => "0000000000000000",
        462 => "0000000000000000",
        463 => "0000000000000000",
        464 => "0000000000000000",
        465 => "0000000000000000",
        466 => "0000000000000000",
        467 => "0000000000000000",
        468 => "0000000000000000",
        469 => "0000000000000000",
        470 => "0000000000000000",
        471 => "0000000000000000",
        472 => "0000000000000000",
        473 => "0000000000000000",
        474 => "0000000000000000",
        475 => "0000000000000000",
        476 => "0000000000000000",
        477 => "0000000000000000",
        478 => "0000000000000000",
        479 => "0000000000000000",
        480 => "0000000000000000",
        481 => "0000000000000000",
        482 => "0000000000000000",
        483 => "0000000000000000",
        484 => "0000000000000000",
        485 => "0000000000000000",
        486 => "0000000000000000",
        487 => "0000000000000000",
        488 => "0000000000000000",
        489 => "0000000000000000",
        490 => "0000000000000000",
        491 => "0000000000000000",
        492 => "0000000000000000",
        493 => "0000000000000000",
        494 => "0000000000000000",
        495 => "0000000000000000",
        496 => "0000000000000000",
        497 => "0000000000000000",
        498 => "0000000000000000",
        499 => "0000000000000000",
        500 => "0000000000000000",
        501 => "0000000000000000",
        502 => "0000000000000000",
        503 => "0000000000000000",
        504 => "0000000000000000",
        505 => "0000000000000000",
        506 => "0000000000000000",
        507 => "0000000000000000",
        508 => "0000000000000000",
        509 => "0000000000000000",
        510 => "0000000000000000",
        511 => "0000000000000000",
        512 => "1000111000000000",
        513 => "1110000011000000",
        514 => "1111000010000000",
        515 => "0010011011000000",
        516 => "0000000000000000",
        517 => "0000000000000000",
        518 => "0000000000000000",
        519 => "0000000000000000",
        520 => "0000000000000000",
        521 => "0000000000000000",
        522 => "0000000000000000",
        523 => "0000000000000000",
        524 => "0000000000000000",
        525 => "0000000000000000",
        526 => "0000000000000000",
        527 => "0000000000000000",
        528 => "0000000000000000",
        529 => "0000000000000000",
        530 => "0000000000000000",
        531 => "0000000000000000",
        532 => "0000000000000000",
        533 => "0000000000000000",
        534 => "0000000000000000",
        535 => "0000000000000000",
        536 => "0000000000000000",
        537 => "0000000000000000",
        538 => "0000000000000000",
        539 => "0000000000000000",
        540 => "0000000000000000",
        541 => "0000000000000000",
        542 => "0000000000000000",
        543 => "0000000000000000",
        544 => "0000000000000000",
        545 => "0000000000000000",
        546 => "0000000000000000",
        547 => "0000000000000000",
        548 => "0000000000000000",
        549 => "0000000000000000",
        550 => "0000000000000000",
        551 => "0000000000000000",
        552 => "0000000000000000",
        553 => "0000000000000000",
        554 => "0000000000000000",
        555 => "0000000000000000",
        556 => "0000000000000000",
        557 => "0000000000000000",
        558 => "0000000000000000",
        559 => "0000000000000000",
        560 => "0000000000000000",
        561 => "0000000000000000",
        562 => "0000000000000000",
        563 => "0000000000000000",
        564 => "0000000000000000",
        565 => "0000000000000000",
        566 => "0000000000000000",
        567 => "0000000000000000",
        568 => "0000000000000000",
        569 => "0000000000000000",
        570 => "0000000000000000",
        571 => "0000000000000000",
        572 => "0000000000000000",
        573 => "0000000000000000",
        574 => "0000000000000000",
        575 => "0000000000000000",
        576 => "0000000000000000",
        577 => "0000000000000000",
        578 => "0000000000000000",
        579 => "0000000000000000",
        580 => "0000000000000000",
        581 => "0000000000000000",
        582 => "0000000000000000",
        583 => "0000000000000000",
        584 => "0000000000000000",
        585 => "0000000000000000",
        586 => "0000000000000000",
        587 => "0000000000000000",
        588 => "0000000000000000",
        589 => "0000000000000000",
        590 => "0000000000000000",
        591 => "0000000000000000",
        592 => "0000000000000000",
        593 => "0000000000000000",
        594 => "0000000000000000",
        595 => "0000000000000000",
        596 => "0000000000000000",
        597 => "0000000000000000",
        598 => "0000000000000000",
        599 => "0000000000000000",
        600 => "0000000000000000",
        601 => "0000000000000000",
        602 => "0000000000000000",
        603 => "0000000000000000",
        604 => "0000000000000000",
        605 => "0000000000000000",
        606 => "0000000000000000",
        607 => "0000000000000000",
        608 => "0000000000000000",
        609 => "0000000000000000",
        610 => "0000000000000000",
        611 => "0000000000000000",
        612 => "0000000000000000",
        613 => "0000000000000000",
        614 => "0000000000000000",
        615 => "0000000000000000",
        616 => "0000000000000000",
        617 => "0000000000000000",
        618 => "0000000000000000",
        619 => "0000000000000000",
        620 => "0000000000000000",
        621 => "0000000000000000",
        622 => "0000000000000000",
        623 => "0000000000000000",
        624 => "0000000000000000",
        625 => "0000000000000000",
        626 => "0000000000000000",
        627 => "0000000000000000",
        628 => "0000000000000000",
        629 => "0000000000000000",
        630 => "0000000000000000",
        631 => "0000000000000000",
        632 => "0000000000000000",
        633 => "0000000000000000",
        634 => "0000000000000000",
        635 => "0000000000000000",
        636 => "0000000000000000",
        637 => "0000000000000000",
        638 => "0000000000000000",
        639 => "0000000000000000",
        640 => "0000000000000000",
        641 => "0000000000000000",
        642 => "0000000000000000",
        643 => "0000000000000000",
        644 => "0000000000000000",
        645 => "0000000000000000",
        646 => "0000000000000000",
        647 => "0000000000000000",
        648 => "0000000000000000",
        649 => "0000000000000000",
        650 => "0000000000000000",
        651 => "0000000000000000",
        652 => "0000000000000000",
        653 => "0000000000000000",
        654 => "0000000000000000",
        655 => "0000000000000000",
        656 => "0000000000000000",
        657 => "0000000000000000",
        658 => "0000000000000000",
        659 => "0000000000000000",
        660 => "0000000000000000",
        661 => "0000000000000000",
        662 => "0000000000000000",
        663 => "0000000000000000",
        664 => "0000000000000000",
        665 => "0000000000000000",
        666 => "0000000000000000",
        667 => "0000000000000000",
        668 => "0000000000000000",
        669 => "0000000000000000",
        670 => "0000000000000000",
        671 => "0000000000000000",
        672 => "0000000000000000",
        673 => "0000000000000000",
        674 => "0000000000000000",
        675 => "0000000000000000",
        676 => "0000000000000000",
        677 => "0000000000000000",
        678 => "0000000000000000",
        679 => "0000000000000000",
        680 => "0000000000000000",
        681 => "0000000000000000",
        682 => "0000000000000000",
        683 => "0000000000000000",
        684 => "0000000000000000",
        685 => "0000000000000000",
        686 => "0000000000000000",
        687 => "0000000000000000",
        688 => "0000000000000000",
        689 => "0000000000000000",
        690 => "0000000000000000",
        691 => "0000000000000000",
        692 => "0000000000000000",
        693 => "0000000000000000",
        694 => "0000000000000000",
        695 => "0000000000000000",
        696 => "0000000000000000",
        697 => "0000000000000000",
        698 => "0000000000000000",
        699 => "0000000000000000",
        700 => "0000000000000000",
        701 => "0000000000000000",
        702 => "0000000000000000",
        703 => "0000000000000000",
        704 => "0000000000000000",
        705 => "0000000000000000",
        706 => "0000000000000000",
        707 => "0000000000000000",
        708 => "0000000000000000",
        709 => "0000000000000000",
        710 => "0000000000000000",
        711 => "0000000000000000",
        712 => "0000000000000000",
        713 => "0000000000000000",
        714 => "0000000000000000",
        715 => "0000000000000000",
        716 => "0000000000000000",
        717 => "0000000000000000",
        718 => "0000000000000000",
        719 => "0000000000000000",
        720 => "0000000000000000",
        721 => "0000000000000000",
        722 => "0000000000000000",
        723 => "0000000000000000",
        724 => "0000000000000000",
        725 => "0000000000000000",
        726 => "0000000000000000",
        727 => "0000000000000000",
        728 => "0000000000000000",
        729 => "0000000000000000",
        730 => "0000000000000000",
        731 => "0000000000000000",
        732 => "0000000000000000",
        733 => "0000000000000000",
        734 => "0000000000000000",
        735 => "0000000000000000",
        736 => "0000000000000000",
        737 => "0000000000000000",
        738 => "0000000000000000",
        739 => "0000000000000000",
        740 => "0000000000000000",
        741 => "0000000000000000",
        742 => "0000000000000000",
        743 => "0000000000000000",
        744 => "0000000000000000",
        745 => "0000000000000000",
        746 => "0000000000000000",
        747 => "0000000000000000",
        748 => "0000000000000000",
        749 => "0000000000000000",
        750 => "0000000000000000",
        751 => "0000000000000000",
        752 => "0000000000000000",
        753 => "0000000000000000",
        754 => "0000000000000000",
        755 => "0000000000000000",
        756 => "0000000000000000",
        757 => "0000000000000000",
        758 => "0000000000000000",
        759 => "0000000000000000",
        760 => "0000000000000000",
        761 => "0000000000000000",
        762 => "0000000000000000",
        763 => "0000000000000000",
        764 => "0000000000000000",
        765 => "0000000000000000",
        766 => "0000000000000000",
        767 => "0000000000000000",
        768 => "0100111001111000",
        769 => "0100100100101000",
        770 => "1110100000000000",
        771 => "0010011111100000",
        772 => "0000000000000000",
        773 => "0000000000000000",
        774 => "0000000000000000",
        775 => "0000000000000000",
        776 => "0000000000000000",
        777 => "0000000000000000",
        778 => "0000000000000000",
        779 => "0000000000000000",
        780 => "0000000000000000",
        781 => "0000000000000000",
        782 => "0000000000000000",
        783 => "0000000000000000",
        784 => "0000000000000000",
        785 => "0000000000000000",
        786 => "0000000000000000",
        787 => "0000000000000000",
        788 => "0000000000000000",
        789 => "0000000000000000",
        790 => "0000000000000000",
        791 => "0000000000000000",
        792 => "0000000000000000",
        793 => "0000000000000000",
        794 => "0000000000000000",
        795 => "0000000000000000",
        796 => "0000000000000000",
        797 => "0000000000000000",
        798 => "0000000000000000",
        799 => "0000000000000000",
        800 => "0000000000000000",
        801 => "0000000000000000",
        802 => "0000000000000000",
        803 => "0000000000000000",
        804 => "0000000000000000",
        805 => "0000000000000000",
        806 => "0000000000000000",
        807 => "0000000000000000",
        808 => "0000000000000000",
        809 => "0000000000000000",
        810 => "0000000000000000",
        811 => "0000000000000000",
        812 => "0000000000000000",
        813 => "0000000000000000",
        814 => "0000000000000000",
        815 => "0000000000000000",
        816 => "0000000000000000",
        817 => "0000000000000000",
        818 => "0000000000000000",
        819 => "0000000000000000",
        820 => "0000000000000000",
        821 => "0000000000000000",
        822 => "0000000000000000",
        823 => "0000000000000000",
        824 => "0000000000000000",
        825 => "0000000000000000",
        826 => "0000000000000000",
        827 => "0000000000000000",
        828 => "0000000000000000",
        829 => "0000000000000000",
        830 => "0000000000000000",
        831 => "0000000000000000",
        832 => "0000000000000000",
        833 => "0000000000000000",
        834 => "0000000000000000",
        835 => "0000000000000000",
        836 => "0000000000000000",
        837 => "0000000000000000",
        838 => "0000000000000000",
        839 => "0000000000000000",
        840 => "0000000000000000",
        841 => "0000000000000000",
        842 => "0000000000000000",
        843 => "0000000000000000",
        844 => "0000000000000000",
        845 => "0000000000000000",
        846 => "0000000000000000",
        847 => "0000000000000000",
        848 => "0000000000000000",
        849 => "0000000000000000",
        850 => "0000000000000000",
        851 => "0000000000000000",
        852 => "0000000000000000",
        853 => "0000000000000000",
        854 => "0000000000000000",
        855 => "0000000000000000",
        856 => "0000000000000000",
        857 => "0000000000000000",
        858 => "0000000000000000",
        859 => "0000000000000000",
        860 => "0000000000000000",
        861 => "0000000000000000",
        862 => "0000000000000000",
        863 => "0000000000000000",
        864 => "0000000000000000",
        865 => "0000000000000000",
        866 => "0000000000000000",
        867 => "0000000000000000",
        868 => "0000000000000000",
        869 => "0000000000000000",
        870 => "0000000000000000",
        871 => "0000000000000000",
        872 => "0000000000000000",
        873 => "0000000000000000",
        874 => "0000000000000000",
        875 => "0000000000000000",
        876 => "0000000000000000",
        877 => "0000000000000000",
        878 => "0000000000000000",
        879 => "0000000000000000",
        880 => "0000000000000000",
        881 => "0000000000000000",
        882 => "0000000000000000",
        883 => "0000000000000000",
        884 => "0000000000000000",
        885 => "0000000000000000",
        886 => "0000000000000000",
        887 => "0000000000000000",
        888 => "0000000000000000",
        889 => "0000000000000000",
        890 => "0000000000000000",
        891 => "0000000000000000",
        892 => "0000000000000000",
        893 => "0000000000000000",
        894 => "0000000000000000",
        895 => "0000000000000000",
        896 => "0000000000000000",
        897 => "0000000000000000",
        898 => "0000000000000000",
        899 => "0000000000000000",
        900 => "0000000000000000",
        901 => "0000000000000000",
        902 => "0000000000000000",
        903 => "0000000000000000",
        904 => "0000000000000000",
        905 => "0000000000000000",
        906 => "0000000000000000",
        907 => "0000000000000000",
        908 => "0000000000000000",
        909 => "0000000000000000",
        910 => "0000000000000000",
        911 => "0000000000000000",
        912 => "0000000000000000",
        913 => "0000000000000000",
        914 => "0000000000000000",
        915 => "0000000000000000",
        916 => "0000000000000000",
        917 => "0000000000000000",
        918 => "0000000000000000",
        919 => "0000000000000000",
        920 => "0000000000000000",
        921 => "0000000000000000",
        922 => "0000000000000000",
        923 => "0000000000000000",
        924 => "0000000000000000",
        925 => "0000000000000000",
        926 => "0000000000000000",
        927 => "0000000000000000",
        928 => "0000000000000000",
        929 => "0000000000000000",
        930 => "0000000000000000",
        931 => "0000000000000000",
        932 => "0000000000000000",
        933 => "0000000000000000",
        934 => "0000000000000000",
        935 => "0000000000000000",
        936 => "0000000000000000",
        937 => "0000000000000000",
        938 => "0000000000000000",
        939 => "0000000000000000",
        940 => "0000000000000000",
        941 => "0000000000000000",
        942 => "0000000000000000",
        943 => "0000000000000000",
        944 => "0000000000000000",
        945 => "0000000000000000",
        946 => "0000000000000000",
        947 => "0000000000000000",
        948 => "0000000000000000",
        949 => "0000000000000000",
        950 => "0000000000000000",
        951 => "0000000000000000",
        952 => "0000000000000000",
        953 => "0000000000000000",
        954 => "0000000000000000",
        955 => "0000000000000000",
        956 => "0000000000000000",
        957 => "0000000000000000",
        958 => "0000000000000000",
        959 => "0000000000000000",
        960 => "0000000000000000",
        961 => "0000000000000000",
        962 => "0000000000000000",
        963 => "0000000000000000",
        964 => "0000000000000000",
        965 => "0000000000000000",
        966 => "0000000000000000",
        967 => "0000000000000000",
        968 => "0000000000000000",
        969 => "0000000000000000",
        970 => "0000000000000000",
        971 => "0000000000000000",
        972 => "0000000000000000",
        973 => "0000000000000000",
        974 => "0000000000000000",
        975 => "0000000000000000",
        976 => "0000000000000000",
        977 => "0000000000000000",
        978 => "0000000000000000",
        979 => "0000000000000000",
        980 => "0000000000000000",
        981 => "0000000000000000",
        982 => "0000000000000000",
        983 => "0000000000000000",
        984 => "0000000000000000",
        985 => "0000000000000000",
        986 => "0000000000000000",
        987 => "0000000000000000",
        988 => "0000000000000000",
        989 => "0000000000000000",
        990 => "0000000000000000",
        991 => "0000000000000000",
        992 => "0000000000000000",
        993 => "0000000000000000",
        994 => "0000000000000000",
        995 => "0000000000000000",
        996 => "0000000000000000",
        997 => "0000000000000000",
        998 => "0000000000000000",
        999 => "0000000000000000",
        1000 => "0000000000000000",
        1001 => "0000000000000000",
        1002 => "0000000000000000",
        1003 => "0000000000000000",
        1004 => "0000000000000000",
        1005 => "0000000000000000",
        1006 => "0000000000000000",
        1007 => "0000000000000000",
        1008 => "0000000000000000",
        1009 => "0000000000000000",
        1010 => "0000000000000000",
        1011 => "0000000000000000",
        1012 => "0000000000000000",
        1013 => "0000000000000000",
        1014 => "0000000000000000",
        1015 => "0000000000000000",
        1016 => "0000000000000000",
        1017 => "0000000000000000",
        1018 => "0000000000000000",
        1019 => "0000000000000000",
        1020 => "0000000000000000",
        1021 => "0000000000000000",
        1022 => "0000000000000000",
        1023 => "0000000000000000",
        1024 => "0000000000000000",
        1025 => "0000100000000000",
        1026 => "0000000000000000",
        1027 => "0000000000000000",
        1028 => "0000000000000000",
        1029 => "0000000000000000",
        1030 => "0000000000000000",
        1031 => "0000000000000000",
        1032 => "0000000000000000",
        1033 => "0000000000000000",
        1034 => "0000000000000000",
        1035 => "0000000000000000",
        1036 => "0000000000000000",
        1037 => "0000000000000000",
        1038 => "0000000000000000",
        1039 => "0000000000000000",
        1040 => "0000000000000000",
        1041 => "0000000000000000",
        1042 => "0000000000000000",
        1043 => "0000000000000000",
        1044 => "0000000000000000",
        1045 => "0000000000000000",
        1046 => "0000000000000000",
        1047 => "0000000000000000",
        1048 => "0000000000000000",
        1049 => "0000000000000000",
        1050 => "0000000000000000",
        1051 => "0000000000000000",
        1052 => "0000000000000000",
        1053 => "0000000000000000",
        1054 => "0000000000000000",
        1055 => "0000000000000000",
        1056 => "0000000000000000",
        1057 => "0000000000000000",
        1058 => "0000000000000000",
        1059 => "0000000000000000",
        1060 => "0000000000000000",
        1061 => "0000000000000000",
        1062 => "0000000000000000",
        1063 => "0000000000000000",
        1064 => "0000000000000000",
        1065 => "0000000000000000",
        1066 => "0000000000000000",
        1067 => "0000000000000000",
        1068 => "0000000000000000",
        1069 => "0000000000000000",
        1070 => "0000000000000000",
        1071 => "0000000000000000",
        1072 => "0000000000000000",
        1073 => "0000000000000000",
        1074 => "0000000000000000",
        1075 => "0000000000000000",
        1076 => "0000000000000000",
        1077 => "0000000000000000",
        1078 => "0000000000000000",
        1079 => "0000000000000000",
        1080 => "0000000000000000",
        1081 => "0000000000000000",
        1082 => "0000000000000000",
        1083 => "0000000000000000",
        1084 => "0000000000000000",
        1085 => "0000000000000000",
        1086 => "0000000000000000",
        1087 => "0000000000000000",
        1088 => "0000000000000000",
        1089 => "0000000000000000",
        1090 => "0000000000000000",
        1091 => "0000000000000000",
        1092 => "0000000000000000",
        1093 => "0000000000000000",
        1094 => "0000000000000000",
        1095 => "0000000000000000",
        1096 => "0000000000000000",
        1097 => "0000000000000000",
        1098 => "0000000000000000",
        1099 => "0000000000000000",
        1100 => "0000000000000000",
        1101 => "0000000000000000",
        1102 => "0000000000000000",
        1103 => "0000000000000000",
        1104 => "0000000000000000",
        1105 => "0000000000000000",
        1106 => "0000000000000000",
        1107 => "0000000000000000",
        1108 => "0000000000000000",
        1109 => "0000000000000000",
        1110 => "0000000000000000",
        1111 => "0000000000000000",
        1112 => "0000000000000000",
        1113 => "0000000000000000",
        1114 => "0000000000000000",
        1115 => "0000000000000000",
        1116 => "0000000000000000",
        1117 => "0000000000000000",
        1118 => "0000000000000000",
        1119 => "0000000000000000",
        1120 => "0000000000000000",
        1121 => "0000000000000000",
        1122 => "0000000000000000",
        1123 => "0000000000000000",
        1124 => "0000000000000000",
        1125 => "0000000000000000",
        1126 => "0000000000000000",
        1127 => "0000000000000000",
        1128 => "0000000000000000",
        1129 => "0000000000000000",
        1130 => "0000000000000000",
        1131 => "0000000000000000",
        1132 => "0000000000000000",
        1133 => "0000000000000000",
        1134 => "0000000000000000",
        1135 => "0000000000000000",
        1136 => "0000000000000000",
        1137 => "0000000000000000",
        1138 => "0000000000000000",
        1139 => "0000000000000000",
        1140 => "0000000000000000",
        1141 => "0000000000000000",
        1142 => "0000000000000000",
        1143 => "0000000000000000",
        1144 => "0000000000000000",
        1145 => "0000000000000000",
        1146 => "0000000000000000",
        1147 => "0000000000000000",
        1148 => "0000000000000000",
        1149 => "0000000000000000",
        1150 => "0000000000000000",
        1151 => "0000000000000000",
        1152 => "0000000000000000",
        1153 => "0000000000000000",
        1154 => "0000000000000000",
        1155 => "0000000000000000",
        1156 => "0000000000000000",
        1157 => "0000000000000000",
        1158 => "0000000000000000",
        1159 => "0000000000000000",
        1160 => "0000000000000000",
        1161 => "0000000000000000",
        1162 => "0000000000000000",
        1163 => "0000000000000000",
        1164 => "0000000000000000",
        1165 => "0000000000000000",
        1166 => "0000000000000000",
        1167 => "0000000000000000",
        1168 => "0000000000000000",
        1169 => "0000000000000000",
        1170 => "0000000000000000",
        1171 => "0000000000000000",
        1172 => "0000000000000000",
        1173 => "0000000000000000",
        1174 => "0000000000000000",
        1175 => "0000000000000000",
        1176 => "0000000000000000",
        1177 => "0000000000000000",
        1178 => "0000000000000000",
        1179 => "0000000000000000",
        1180 => "0000000000000000",
        1181 => "0000000000000000",
        1182 => "0000000000000000",
        1183 => "0000000000000000",
        1184 => "0000000000000000",
        1185 => "0000000000000000",
        1186 => "0000000000000000",
        1187 => "0000000000000000",
        1188 => "0000000000000000",
        1189 => "0000000000000000",
        1190 => "0000000000000000",
        1191 => "0000000000000000",
        1192 => "0000000000000000",
        1193 => "0000000000000000",
        1194 => "0000000000000000",
        1195 => "0000000000000000",
        1196 => "0000000000000000",
        1197 => "0000000000000000",
        1198 => "0000000000000000",
        1199 => "0000000000000000",
        1200 => "0000000000000000",
        1201 => "0000000000000000",
        1202 => "0000000000000000",
        1203 => "0000000000000000",
        1204 => "0000000000000000",
        1205 => "0000000000000000",
        1206 => "0000000000000000",
        1207 => "0000000000000000",
        1208 => "0000000000000000",
        1209 => "0000000000000000",
        1210 => "0000000000000000",
        1211 => "0000000000000000",
        1212 => "0000000000000000",
        1213 => "0000000000000000",
        1214 => "0000000000000000",
        1215 => "0000000000000000",
        1216 => "0000000000000000",
        1217 => "0000000000000000",
        1218 => "0000000000000000",
        1219 => "0000000000000000",
        1220 => "0000000000000000",
        1221 => "0000000000000000",
        1222 => "0000000000000000",
        1223 => "0000000000000000",
        1224 => "0000000000000000",
        1225 => "0000000000000000",
        1226 => "0000000000000000",
        1227 => "0000000000000000",
        1228 => "0000000000000000",
        1229 => "0000000000000000",
        1230 => "0000000000000000",
        1231 => "0000000000000000",
        1232 => "0000000000000000",
        1233 => "0000000000000000",
        1234 => "0000000000000000",
        1235 => "0000000000000000",
        1236 => "0000000000000000",
        1237 => "0000000000000000",
        1238 => "0000000000000000",
        1239 => "0000000000000000",
        1240 => "0000000000000000",
        1241 => "0000000000000000",
        1242 => "0000000000000000",
        1243 => "0000000000000000",
        1244 => "0000000000000000",
        1245 => "0000000000000000",
        1246 => "0000000000000000",
        1247 => "0000000000000000",
        1248 => "0000000000000000",
        1249 => "0000000000000000",
        1250 => "0000000000000000",
        1251 => "0000000000000000",
        1252 => "0000000000000000",
        1253 => "0000000000000000",
        1254 => "0000000000000000",
        1255 => "0000000000000000",
        1256 => "0000000000000000",
        1257 => "0000000000000000",
        1258 => "0000000000000000",
        1259 => "0000000000000000",
        1260 => "0000000000000000",
        1261 => "0000000000000000",
        1262 => "0000000000000000",
        1263 => "0000000000000000",
        1264 => "0000000000000000",
        1265 => "0000000000000000",
        1266 => "0000000000000000",
        1267 => "0000000000000000",
        1268 => "0000000000000000",
        1269 => "0000000000000000",
        1270 => "0000000000000000",
        1271 => "0000000000000000",
        1272 => "0000000000000000",
        1273 => "0000000000000000",
        1274 => "0000000000000000",
        1275 => "0000000000000000",
        1276 => "0000000000000000",
        1277 => "0000000000000000",
        1278 => "0000000000000000",
        1279 => "0000000000000000",
        1280 => "0000000000000000",
        1281 => "0000000000000000",
        1282 => "0000000000000000",
        1283 => "0000000000000000",
        1284 => "0000000000000000",
        1285 => "0000000000000000",
        1286 => "0000000000000000",
        1287 => "0000000000000000",
        1288 => "0000000000000000",
        1289 => "0000000000000000",
        1290 => "0000000000000000",
        1291 => "0000000000000000",
        1292 => "0000000000000000",
        1293 => "0000000000000000",
        1294 => "0000000000000000",
        1295 => "0000000000000000",
        1296 => "0000000000000000",
        1297 => "0000000000000000",
        1298 => "0000000000000000",
        1299 => "0000000000000000",
        1300 => "0000000000000000",
        1301 => "0000000000000000",
        1302 => "0000000000000000",
        1303 => "0000000000000000",
        1304 => "0000000000000000",
        1305 => "0000000000000000",
        1306 => "0000000000000000",
        1307 => "0000000000000000",
        1308 => "0000000000000000",
        1309 => "0000000000000000",
        1310 => "0000000000000000",
        1311 => "0000000000000000",
        1312 => "0000000000000000",
        1313 => "0000000000000000",
        1314 => "0000000000000000",
        1315 => "0000000000000000",
        1316 => "0000000000000000",
        1317 => "0000000000000000",
        1318 => "0000000000000000",
        1319 => "0000000000000000",
        1320 => "0000000000000000",
        1321 => "0000000000000000",
        1322 => "0000000000000000",
        1323 => "0000000000000000",
        1324 => "0000000000000000",
        1325 => "0000000000000000",
        1326 => "0000000000000000",
        1327 => "0000000000000000",
        1328 => "0000000000000000",
        1329 => "0000000000000000",
        1330 => "0000000000000000",
        1331 => "0000000000000000",
        1332 => "0000000000000000",
        1333 => "0000000000000000",
        1334 => "0000000000000000",
        1335 => "0000000000000000",
        1336 => "0000000000000000",
        1337 => "0000000000000000",
        1338 => "0000000000000000",
        1339 => "0000000000000000",
        1340 => "0000000000000000",
        1341 => "0000000000000000",
        1342 => "0000000000000000",
        1343 => "0000000000000000",
        1344 => "0000000000000000",
        1345 => "0000000000000000",
        1346 => "0000000000000000",
        1347 => "0000000000000000",
        1348 => "0000000000000000",
        1349 => "0000000000000000",
        1350 => "0000000000000000",
        1351 => "0000000000000000",
        1352 => "0000000000000000",
        1353 => "0000000000000000",
        1354 => "0000000000000000",
        1355 => "0000000000000000",
        1356 => "0000000000000000",
        1357 => "0000000000000000",
        1358 => "0000000000000000",
        1359 => "0000000000000000",
        1360 => "0000000000000000",
        1361 => "0000000000000000",
        1362 => "0000000000000000",
        1363 => "0000000000000000",
        1364 => "0000000000000000",
        1365 => "0000000000000000",
        1366 => "0000000000000000",
        1367 => "0000000000000000",
        1368 => "0000000000000000",
        1369 => "0000000000000000",
        1370 => "0000000000000000",
        1371 => "0000000000000000",
        1372 => "0000000000000000",
        1373 => "0000000000000000",
        1374 => "0000000000000000",
        1375 => "0000000000000000",
        1376 => "0000000000000000",
        1377 => "0000000000000000",
        1378 => "0000000000000000",
        1379 => "0000000000000000",
        1380 => "0000000000000000",
        1381 => "0000000000000000",
        1382 => "0000000000000000",
        1383 => "0000000000000000",
        1384 => "0000000000000000",
        1385 => "0000000000000000",
        1386 => "0000000000000000",
        1387 => "0000000000000000",
        1388 => "0000000000000000",
        1389 => "0000000000000000",
        1390 => "0000000000000000",
        1391 => "0000000000000000",
        1392 => "0000000000000000",
        1393 => "0000000000000000",
        1394 => "0000000000000000",
        1395 => "0000000000000000",
        1396 => "0000000000000000",
        1397 => "0000000000000000",
        1398 => "0000000000000000",
        1399 => "0000000000000000",
        1400 => "0000000000000000",
        1401 => "0000000000000000",
        1402 => "0000000000000000",
        1403 => "0000000000000000",
        1404 => "0000000000000000",
        1405 => "0000000000000000",
        1406 => "0000000000000000",
        1407 => "0000000000000000",
        1408 => "0000000000000000",
        1409 => "0000000000000000",
        1410 => "0000000000000000",
        1411 => "0000000000000000",
        1412 => "0000000000000000",
        1413 => "0000000000000000",
        1414 => "0000000000000000",
        1415 => "0000000000000000",
        1416 => "0000000000000000",
        1417 => "0000000000000000",
        1418 => "0000000000000000",
        1419 => "0000000000000000",
        1420 => "0000000000000000",
        1421 => "0000000000000000",
        1422 => "0000000000000000",
        1423 => "0000000000000000",
        1424 => "0000000000000000",
        1425 => "0000000000000000",
        1426 => "0000000000000000",
        1427 => "0000000000000000",
        1428 => "0000000000000000",
        1429 => "0000000000000000",
        1430 => "0000000000000000",
        1431 => "0000000000000000",
        1432 => "0000000000000000",
        1433 => "0000000000000000",
        1434 => "0000000000000000",
        1435 => "0000000000000000",
        1436 => "0000000000000000",
        1437 => "0000000000000000",
        1438 => "0000000000000000",
        1439 => "0000000000000000",
        1440 => "0000000000000000",
        1441 => "0000000000000000",
        1442 => "0000000000000000",
        1443 => "0000000000000000",
        1444 => "0000000000000000",
        1445 => "0000000000000000",
        1446 => "0000000000000000",
        1447 => "0000000000000000",
        1448 => "0000000000000000",
        1449 => "0000000000000000",
        1450 => "0000000000000000",
        1451 => "0000000000000000",
        1452 => "0000000000000000",
        1453 => "0000000000000000",
        1454 => "0000000000000000",
        1455 => "0000000000000000",
        1456 => "0000000000000000",
        1457 => "0000000000000000",
        1458 => "0000000000000000",
        1459 => "0000000000000000",
        1460 => "0000000000000000",
        1461 => "0000000000000000",
        1462 => "0000000000000000",
        1463 => "0000000000000000",
        1464 => "0000000000000000",
        1465 => "0000000000000000",
        1466 => "0000000000000000",
        1467 => "0000000000000000",
        1468 => "0000000000000000",
        1469 => "0000000000000000",
        1470 => "0000000000000000",
        1471 => "0000000000000000",
        1472 => "0000000000000000",
        1473 => "0000000000000000",
        1474 => "0000000000000000",
        1475 => "0000000000000000",
        1476 => "0000000000000000",
        1477 => "0000000000000000",
        1478 => "0000000000000000",
        1479 => "0000000000000000",
        1480 => "0000000000000000",
        1481 => "0000000000000000",
        1482 => "0000000000000000",
        1483 => "0000000000000000",
        1484 => "0000000000000000",
        1485 => "0000000000000000",
        1486 => "0000000000000000",
        1487 => "0000000000000000",
        1488 => "0000000000000000",
        1489 => "0000000000000000",
        1490 => "0000000000000000",
        1491 => "0000000000000000",
        1492 => "0000000000000000",
        1493 => "0000000000000000",
        1494 => "0000000000000000",
        1495 => "0000000000000000",
        1496 => "0000000000000000",
        1497 => "0000000000000000",
        1498 => "0000000000000000",
        1499 => "0000000000000000",
        1500 => "0000000000000000",
        1501 => "0000000000000000",
        1502 => "0000000000000000",
        1503 => "0000000000000000",
        1504 => "0000000000000000",
        1505 => "0000000000000000",
        1506 => "0000000000000000",
        1507 => "0000000000000000",
        1508 => "0000000000000000",
        1509 => "0000000000000000",
        1510 => "0000000000000000",
        1511 => "0000000000000000",
        1512 => "0000000000000000",
        1513 => "0000000000000000",
        1514 => "0000000000000000",
        1515 => "0000000000000000",
        1516 => "0000000000000000",
        1517 => "0000000000000000",
        1518 => "0000000000000000",
        1519 => "0000000000000000",
        1520 => "0000000000000000",
        1521 => "0000000000000000",
        1522 => "0000000000000000",
        1523 => "0000000000000000",
        1524 => "0000000000000000",
        1525 => "0000000000000000",
        1526 => "0000000000000000",
        1527 => "0000000000000000",
        1528 => "0000000000000000",
        1529 => "0000000000000000",
        1530 => "0000000000000000",
        1531 => "0000000000000000",
        1532 => "0000000000000000",
        1533 => "0000000000000000",
        1534 => "0000000000000000",
        1535 => "0000000000000000",
        1536 => "0000000000000000",
        1537 => "0000100000000000",
        1538 => "0000000000000000",
        1539 => "0000000000000000",
        1540 => "0000000000000000",
        1541 => "0000000000000000",
        1542 => "0000000000000000",
        1543 => "0000000000000000",
        1544 => "0000000000000000",
        1545 => "0000000000000000",
        1546 => "0000000000000000",
        1547 => "0000000000000000",
        1548 => "0000000000000000",
        1549 => "0000000000000000",
        1550 => "0000000000000000",
        1551 => "0000000000000000",
        1552 => "0000000000000000",
        1553 => "0000000000000000",
        1554 => "0000000000000000",
        1555 => "0000000000000000",
        1556 => "0000000000000000",
        1557 => "0000000000000000",
        1558 => "0000000000000000",
        1559 => "0000000000000000",
        1560 => "0000000000000000",
        1561 => "0000000000000000",
        1562 => "0000000000000000",
        1563 => "0000000000000000",
        1564 => "0000000000000000",
        1565 => "0000000000000000",
        1566 => "0000000000000000",
        1567 => "0000000000000000",
        1568 => "0000000000000000",
        1569 => "0000000000000000",
        1570 => "0000000000000000",
        1571 => "0000000000000000",
        1572 => "0000000000000000",
        1573 => "0000000000000000",
        1574 => "0000000000000000",
        1575 => "0000000000000000",
        1576 => "0000000000000000",
        1577 => "0000000000000000",
        1578 => "0000000000000000",
        1579 => "0000000000000000",
        1580 => "0000000000000000",
        1581 => "0000000000000000",
        1582 => "0000000000000000",
        1583 => "0000000000000000",
        1584 => "0000000000000000",
        1585 => "0000000000000000",
        1586 => "0000000000000000",
        1587 => "0000000000000000",
        1588 => "0000000000000000",
        1589 => "0000000000000000",
        1590 => "0000000000000000",
        1591 => "0000000000000000",
        1592 => "0000000000000000",
        1593 => "0000000000000000",
        1594 => "0000000000000000",
        1595 => "0000000000000000",
        1596 => "0000000000000000",
        1597 => "0000000000000000",
        1598 => "0000000000000000",
        1599 => "0000000000000000",
        1600 => "0000000000000000",
        1601 => "0000000000000000",
        1602 => "0000000000000000",
        1603 => "0000000000000000",
        1604 => "0000000000000000",
        1605 => "0000000000000000",
        1606 => "0000000000000000",
        1607 => "0000000000000000",
        1608 => "0000000000000000",
        1609 => "0000000000000000",
        1610 => "0000000000000000",
        1611 => "0000000000000000",
        1612 => "0000000000000000",
        1613 => "0000000000000000",
        1614 => "0000000000000000",
        1615 => "0000000000000000",
        1616 => "0000000000000000",
        1617 => "0000000000000000",
        1618 => "0000000000000000",
        1619 => "0000000000000000",
        1620 => "0000000000000000",
        1621 => "0000000000000000",
        1622 => "0000000000000000",
        1623 => "0000000000000000",
        1624 => "0000000000000000",
        1625 => "0000000000000000",
        1626 => "0000000000000000",
        1627 => "0000000000000000",
        1628 => "0000000000000000",
        1629 => "0000000000000000",
        1630 => "0000000000000000",
        1631 => "0000000000000000",
        1632 => "0000000000000000",
        1633 => "0000000000000000",
        1634 => "0000000000000000",
        1635 => "0000000000000000",
        1636 => "0000000000000000",
        1637 => "0000000000000000",
        1638 => "0000000000000000",
        1639 => "0000000000000000",
        1640 => "0000000000000000",
        1641 => "0000000000000000",
        1642 => "0000000000000000",
        1643 => "0000000000000000",
        1644 => "0000000000000000",
        1645 => "0000000000000000",
        1646 => "0000000000000000",
        1647 => "0000000000000000",
        1648 => "0000000000000000",
        1649 => "0000000000000000",
        1650 => "0000000000000000",
        1651 => "0000000000000000",
        1652 => "0000000000000000",
        1653 => "0000000000000000",
        1654 => "0000000000000000",
        1655 => "0000000000000000",
        1656 => "0000000000000000",
        1657 => "0000000000000000",
        1658 => "0000000000000000",
        1659 => "0000000000000000",
        1660 => "0000000000000000",
        1661 => "0000000000000000",
        1662 => "0000000000000000",
        1663 => "0000000000000000",
        1664 => "0000000000000000",
        1665 => "0000000000000000",
        1666 => "0000000000000000",
        1667 => "0000000000000000",
        1668 => "0000000000000000",
        1669 => "0000000000000000",
        1670 => "0000000000000000",
        1671 => "0000000000000000",
        1672 => "0000000000000000",
        1673 => "0000000000000000",
        1674 => "0000000000000000",
        1675 => "0000000000000000",
        1676 => "0000000000000000",
        1677 => "0000000000000000",
        1678 => "0000000000000000",
        1679 => "0000000000000000",
        1680 => "0000000000000000",
        1681 => "0000000000000000",
        1682 => "0000000000000000",
        1683 => "0000000000000000",
        1684 => "0000000000000000",
        1685 => "0000000000000000",
        1686 => "0000000000000000",
        1687 => "0000000000000000",
        1688 => "0000000000000000",
        1689 => "0000000000000000",
        1690 => "0000000000000000",
        1691 => "0000000000000000",
        1692 => "0000000000000000",
        1693 => "0000000000000000",
        1694 => "0000000000000000",
        1695 => "0000000000000000",
        1696 => "0000000000000000",
        1697 => "0000000000000000",
        1698 => "0000000000000000",
        1699 => "0000000000000000",
        1700 => "0000000000000000",
        1701 => "0000000000000000",
        1702 => "0000000000000000",
        1703 => "0000000000000000",
        1704 => "0000000000000000",
        1705 => "0000000000000000",
        1706 => "0000000000000000",
        1707 => "0000000000000000",
        1708 => "0000000000000000",
        1709 => "0000000000000000",
        1710 => "0000000000000000",
        1711 => "0000000000000000",
        1712 => "0000000000000000",
        1713 => "0000000000000000",
        1714 => "0000000000000000",
        1715 => "0000000000000000",
        1716 => "0000000000000000",
        1717 => "0000000000000000",
        1718 => "0000000000000000",
        1719 => "0000000000000000",
        1720 => "0000000000000000",
        1721 => "0000000000000000",
        1722 => "0000000000000000",
        1723 => "0000000000000000",
        1724 => "0000000000000000",
        1725 => "0000000000000000",
        1726 => "0000000000000000",
        1727 => "0000000000000000",
        1728 => "0000000000000000",
        1729 => "0000000000000000",
        1730 => "0000000000000000",
        1731 => "0000000000000000",
        1732 => "0000000000000000",
        1733 => "0000000000000000",
        1734 => "0000000000000000",
        1735 => "0000000000000000",
        1736 => "0000000000000000",
        1737 => "0000000000000000",
        1738 => "0000000000000000",
        1739 => "0000000000000000",
        1740 => "0000000000000000",
        1741 => "0000000000000000",
        1742 => "0000000000000000",
        1743 => "0000000000000000",
        1744 => "0000000000000000",
        1745 => "0000000000000000",
        1746 => "0000000000000000",
        1747 => "0000000000000000",
        1748 => "0000000000000000",
        1749 => "0000000000000000",
        1750 => "0000000000000000",
        1751 => "0000000000000000",
        1752 => "0000000000000000",
        1753 => "0000000000000000",
        1754 => "0000000000000000",
        1755 => "0000000000000000",
        1756 => "0000000000000000",
        1757 => "0000000000000000",
        1758 => "0000000000000000",
        1759 => "0000000000000000",
        1760 => "0000000000000000",
        1761 => "0000000000000000",
        1762 => "0000000000000000",
        1763 => "0000000000000000",
        1764 => "0000000000000000",
        1765 => "0000000000000000",
        1766 => "0000000000000000",
        1767 => "0000000000000000",
        1768 => "0000000000000000",
        1769 => "0000000000000000",
        1770 => "0000000000000000",
        1771 => "0000000000000000",
        1772 => "0000000000000000",
        1773 => "0000000000000000",
        1774 => "0000000000000000",
        1775 => "0000000000000000",
        1776 => "0000000000000000",
        1777 => "0000000000000000",
        1778 => "0000000000000000",
        1779 => "0000000000000000",
        1780 => "0000000000000000",
        1781 => "0000000000000000",
        1782 => "0000000000000000",
        1783 => "0000000000000000",
        1784 => "0000000000000000",
        1785 => "0000000000000000",
        1786 => "0000000000000000",
        1787 => "0000000000000000",
        1788 => "0000000000000000",
        1789 => "0000000000000000",
        1790 => "0000000000000000",
        1791 => "0000000000000000",
        1792 => "0011000100000000",
        1793 => "0011001000000000",
        1794 => "0011001100000000",
        1795 => "0011010000000000",
        1796 => "0011011000000000",
        1797 => "0011011100000000",
        1798 => "1000000010000000",
        1799 => "1101100000100000",
        1800 => "0010011111100000",
        1801 => "0000000000000000",
        1802 => "0000000000000000",
        1803 => "0000000000000000",
        1804 => "0000000000000000",
        1805 => "0000000000000000",
        1806 => "0000000000000000",
        1807 => "0000000000000000",
        1808 => "0000000000000000",
        1809 => "0000000000000000",
        1810 => "0000000000000000",
        1811 => "0000000000000000",
        1812 => "0000000000000000",
        1813 => "0000000000000000",
        1814 => "0000000000000000",
        1815 => "0000000000000000",
        1816 => "0000000000000000",
        1817 => "0000000000000000",
        1818 => "0000000000000000",
        1819 => "0000000000000000",
        1820 => "0000000000000000",
        1821 => "0000000000000000",
        1822 => "0000000000000000",
        1823 => "0000000000000000",
        1824 => "0000000000000000",
        1825 => "0000000000000000",
        1826 => "0000000000000000",
        1827 => "0000000000000000",
        1828 => "0000000000000000",
        1829 => "0000000000000000",
        1830 => "0000000000000000",
        1831 => "0000000000000000",
        1832 => "0000000000000000",
        1833 => "0000000000000000",
        1834 => "0000000000000000",
        1835 => "0000000000000000",
        1836 => "0000000000000000",
        1837 => "0000000000000000",
        1838 => "0000000000000000",
        1839 => "0000000000000000",
        1840 => "0000000000000000",
        1841 => "0000000000000000",
        1842 => "0000000000000000",
        1843 => "0000000000000000",
        1844 => "0000000000000000",
        1845 => "0000000000000000",
        1846 => "0000000000000000",
        1847 => "0000000000000000",
        1848 => "0000000000000000",
        1849 => "0000000000000000",
        1850 => "0000000000000000",
        1851 => "0000000000000000",
        1852 => "0000000000000000",
        1853 => "0000000000000000",
        1854 => "0000000000000000",
        1855 => "0000000000000000",
        1856 => "0000000000000000",
        1857 => "0000000000000000",
        1858 => "0000000000000000",
        1859 => "0000000000000000",
        1860 => "0000000000000000",
        1861 => "0000000000000000",
        1862 => "0000000000000000",
        1863 => "0000000000000000",
        1864 => "0000000000000000",
        1865 => "0000000000000000",
        1866 => "0000000000000000",
        1867 => "0000000000000000",
        1868 => "0000000000000000",
        1869 => "0000000000000000",
        1870 => "0000000000000000",
        1871 => "0000000000000000",
        1872 => "0000000000000000",
        1873 => "0000000000000000",
        1874 => "0000000000000000",
        1875 => "0000000000000000",
        1876 => "0000000000000000",
        1877 => "0000000000000000",
        1878 => "0000000000000000",
        1879 => "0000000000000000",
        1880 => "0000000000000000",
        1881 => "0000000000000000",
        1882 => "0000000000000000",
        1883 => "0000000000000000",
        1884 => "0000000000000000",
        1885 => "0000000000000000",
        1886 => "0000000000000000",
        1887 => "0000000000000000",
        1888 => "0000000000000000",
        1889 => "0000000000000000",
        1890 => "0000000000000000",
        1891 => "0000000000000000",
        1892 => "0000000000000000",
        1893 => "0000000000000000",
        1894 => "0000000000000000",
        1895 => "0000000000000000",
        1896 => "0000000000000000",
        1897 => "0000000000000000",
        1898 => "0000000000000000",
        1899 => "0000000000000000",
        1900 => "0000000000000000",
        1901 => "0000000000000000",
        1902 => "0000000000000000",
        1903 => "0000000000000000",
        1904 => "0000000000000000",
        1905 => "0000000000000000",
        1906 => "0000000000000000",
        1907 => "0000000000000000",
        1908 => "0000000000000000",
        1909 => "0000000000000000",
        1910 => "0000000000000000",
        1911 => "0000000000000000",
        1912 => "0000000000000000",
        1913 => "0000000000000000",
        1914 => "0000000000000000",
        1915 => "0000000000000000",
        1916 => "0000000000000000",
        1917 => "0000000000000000",
        1918 => "0000000000000000",
        1919 => "0000000000000000",
        1920 => "0000000000000000",
        1921 => "0000000000000000",
        1922 => "0000000000000000",
        1923 => "0000000000000000",
        1924 => "0000000000000000",
        1925 => "0000000000000000",
        1926 => "0000000000000000",
        1927 => "0000000000000000",
        1928 => "0000000000000000",
        1929 => "0000000000000000",
        1930 => "0000000000000000",
        1931 => "0000000000000000",
        1932 => "0000000000000000",
        1933 => "0000000000000000",
        1934 => "0000000000000000",
        1935 => "0000000000000000",
        1936 => "0000000000000000",
        1937 => "0000000000000000",
        1938 => "0000000000000000",
        1939 => "0000000000000000",
        1940 => "0000000000000000",
        1941 => "0000000000000000",
        1942 => "0000000000000000",
        1943 => "0000000000000000",
        1944 => "0000000000000000",
        1945 => "0000000000000000",
        1946 => "0000000000000000",
        1947 => "0000000000000000",
        1948 => "0000000000000000",
        1949 => "0000000000000000",
        1950 => "0000000000000000",
        1951 => "0000000000000000",
        1952 => "0000000000000000",
        1953 => "0000000000000000",
        1954 => "0000000000000000",
        1955 => "0000000000000000",
        1956 => "0000000000000000",
        1957 => "0000000000000000",
        1958 => "0000000000000000",
        1959 => "0000000000000000",
        1960 => "0000000000000000",
        1961 => "0000000000000000",
        1962 => "0000000000000000",
        1963 => "0000000000000000",
        1964 => "0000000000000000",
        1965 => "0000000000000000",
        1966 => "0000000000000000",
        1967 => "0000000000000000",
        1968 => "0000000000000000",
        1969 => "0000000000000000",
        1970 => "0000000000000000",
        1971 => "0000000000000000",
        1972 => "0000000000000000",
        1973 => "0000000000000000",
        1974 => "0000000000000000",
        1975 => "0000000000000000",
        1976 => "0000000000000000",
        1977 => "0000000000000000",
        1978 => "0000000000000000",
        1979 => "0000000000000000",
        1980 => "0000000000000000",
        1981 => "0000000000000000",
        1982 => "0000000000000000",
        1983 => "0000000000000000",
        1984 => "0000000000000000",
        1985 => "0000000000000000",
        1986 => "0000000000000000",
        1987 => "0000000000000000",
        1988 => "0000000000000000",
        1989 => "0000000000000000",
        1990 => "0000000000000000",
        1991 => "0000000000000000",
        1992 => "0000000000000000",
        1993 => "0000000000000000",
        1994 => "0000000000000000",
        1995 => "0000000000000000",
        1996 => "0000000000000000",
        1997 => "0000000000000000",
        1998 => "0000000000000000",
        1999 => "0000000000000000",
        2000 => "0000000000000000",
        2001 => "0000000000000000",
        2002 => "0000000000000000",
        2003 => "0000000000000000",
        2004 => "0000000000000000",
        2005 => "0000000000000000",
        2006 => "0000000000000000",
        2007 => "0000000000000000",
        2008 => "0000000000000000",
        2009 => "0000000000000000",
        2010 => "0000000000000000",
        2011 => "0000000000000000",
        2012 => "0000000000000000",
        2013 => "0000000000000000",
        2014 => "0000000000000000",
        2015 => "0000000000000000",
        2016 => "0000000000000000",
        2017 => "0000000000000000",
        2018 => "0000000000000000",
        2019 => "0000000000000000",
        2020 => "0000000000000000",
        2021 => "0000000000000000",
        2022 => "0000000000000000",
        2023 => "0000000000000000",
        2024 => "0000000000000000",
        2025 => "0000000000000000",
        2026 => "0000000000000000",
        2027 => "0000000000000000",
        2028 => "0000000000000000",
        2029 => "0000000000000000",
        2030 => "0000000000000000",
        2031 => "0000000000000000",
        2032 => "0000000000000000",
        2033 => "0000000000000000",
        2034 => "0000000000000000",
        2035 => "0000000000000000",
        2036 => "0000000000000000",
        2037 => "0000000000000000",
        2038 => "0000000000000000",
        2039 => "0000000000000000",
        2040 => "0000000000000000",
        2041 => "0000000000000000",
        2042 => "0000000000000000",
        2043 => "0000000000000000",
        2044 => "0000000000000000",
        2045 => "0000000000000000",
        2046 => "0000000000000000",
        2047 => "0000000000000000",
        2048 => "0100100000000000",
        2049 => "0010100011000000",
        2050 => "1111100000000000",
        2051 => "0000000000000000",
        2052 => "0000000000000000",
        2053 => "0000000000000000",
        2054 => "0000000000000000",
        2055 => "0000000000000000",
        2056 => "0000000000000000",
        2057 => "0000000000000000",
        2058 => "0000000000000000",
        2059 => "0000000000000000",
        2060 => "0000000000000000",
        2061 => "0000000000000000",
        2062 => "0000000000000000",
        2063 => "0000000000000000",
        2064 => "0000000000000000",
        2065 => "0000000000000000",
        2066 => "0000000000000000",
        2067 => "0000000000000000",
        2068 => "0000000000000000",
        2069 => "0000000000000000",
        2070 => "0000000000000000",
        2071 => "0000000000000000",
        2072 => "0000000000000000",
        2073 => "0000000000000000",
        2074 => "0000000000000000",
        2075 => "0000000000000000",
        2076 => "0000000000000000",
        2077 => "0000000000000000",
        2078 => "0000000000000000",
        2079 => "0000000000000000",
        2080 => "0000000000000000",
        2081 => "0000000000000000",
        2082 => "0000000000000000",
        2083 => "0000000000000000",
        2084 => "0000000000000000",
        2085 => "0000000000000000",
        2086 => "0000000000000000",
        2087 => "0000000000000000",
        2088 => "0000000000000000",
        2089 => "0000000000000000",
        2090 => "0000000000000000",
        2091 => "0000000000000000",
        2092 => "0000000000000000",
        2093 => "0000000000000000",
        2094 => "0000000000000000",
        2095 => "0000000000000000",
        2096 => "0000000000000000",
        2097 => "0000000000000000",
        2098 => "0000000000000000",
        2099 => "0000000000000000",
        2100 => "0000000000000000",
        2101 => "0000000000000000",
        2102 => "0000000000000000",
        2103 => "0000000000000000",
        2104 => "0000000000000000",
        2105 => "0000000000000000",
        2106 => "0000000000000000",
        2107 => "0000000000000000",
        2108 => "0000000000000000",
        2109 => "0000000000000000",
        2110 => "0000000000000000",
        2111 => "0000000000000000",
        2112 => "0000000000000000",
        2113 => "0000000000000000",
        2114 => "0000000000000000",
        2115 => "0000000000000000",
        2116 => "0000000000000000",
        2117 => "0000000000000000",
        2118 => "0000000000000000",
        2119 => "0000000000000000",
        2120 => "0000000000000000",
        2121 => "0000000000000000",
        2122 => "0000000000000000",
        2123 => "0000000000000000",
        2124 => "0000000000000000",
        2125 => "0000000000000000",
        2126 => "0000000000000000",
        2127 => "0000000000000000",
        2128 => "0000000000000000",
        2129 => "0000000000000000",
        2130 => "0000000000000000",
        2131 => "0000000000000000",
        2132 => "0000000000000000",
        2133 => "0000000000000000",
        2134 => "0000000000000000",
        2135 => "0000000000000000",
        2136 => "0000000000000000",
        2137 => "0000000000000000",
        2138 => "0000000000000000",
        2139 => "0000000000000000",
        2140 => "0000000000000000",
        2141 => "0000000000000000",
        2142 => "0000000000000000",
        2143 => "0000000000000000",
        2144 => "0000000000000000",
        2145 => "0000000000000000",
        2146 => "0000000000000000",
        2147 => "0000000000000000",
        2148 => "0000000000000000",
        2149 => "0000000000000000",
        2150 => "0000000000000000",
        2151 => "0000000000000000",
        2152 => "0000000000000000",
        2153 => "0000000000000000",
        2154 => "0000000000000000",
        2155 => "0000000000000000",
        2156 => "0000000000000000",
        2157 => "0000000000000000",
        2158 => "0000000000000000",
        2159 => "0000000000000000",
        2160 => "0000000000000000",
        2161 => "0000000000000000",
        2162 => "0000000000000000",
        2163 => "0000000000000000",
        2164 => "0000000000000000",
        2165 => "0000000000000000",
        2166 => "0000000000000000",
        2167 => "0000000000000000",
        2168 => "0000000000000000",
        2169 => "0000000000000000",
        2170 => "0000000000000000",
        2171 => "0000000000000000",
        2172 => "0000000000000000",
        2173 => "0000000000000000",
        2174 => "0000000000000000",
        2175 => "0000000000000000",
        2176 => "0000000000000000",
        2177 => "0000000000000000",
        2178 => "0000000000000000",
        2179 => "0000000000000000",
        2180 => "0000000000000000",
        2181 => "0000000000000000",
        2182 => "0000000000000000",
        2183 => "0000000000000000",
        2184 => "0000000000000000",
        2185 => "0000000000000000",
        2186 => "0000000000000000",
        2187 => "0000000000000000",
        2188 => "0000000000000000",
        2189 => "0000000000000000",
        2190 => "0000000000000000",
        2191 => "0000000000000000",
        2192 => "0000000000000000",
        2193 => "0000000000000000",
        2194 => "0000000000000000",
        2195 => "0000000000000000",
        2196 => "0000000000000000",
        2197 => "0000000000000000",
        2198 => "0000000000000000",
        2199 => "0000000000000000",
        2200 => "0000000000000000",
        2201 => "0000000000000000",
        2202 => "0000000000000000",
        2203 => "0000000000000000",
        2204 => "0000000000000000",
        2205 => "0000000000000000",
        2206 => "0000000000000000",
        2207 => "0000000000000000",
        2208 => "0000000000000000",
        2209 => "0000000000000000",
        2210 => "0000000000000000",
        2211 => "0000000000000000",
        2212 => "0000000000000000",
        2213 => "0000000000000000",
        2214 => "0000000000000000",
        2215 => "0000000000000000",
        2216 => "0000000000000000",
        2217 => "0000000000000000",
        2218 => "0000000000000000",
        2219 => "0000000000000000",
        2220 => "0000000000000000",
        2221 => "0000000000000000",
        2222 => "0000000000000000",
        2223 => "0000000000000000",
        2224 => "0000000000000000",
        2225 => "0000000000000000",
        2226 => "0000000000000000",
        2227 => "0000000000000000",
        2228 => "0000000000000000",
        2229 => "0000000000000000",
        2230 => "0000000000000000",
        2231 => "0000000000000000",
        2232 => "0000000000000000",
        2233 => "0000000000000000",
        2234 => "0000000000000000",
        2235 => "0000000000000000",
        2236 => "0000000000000000",
        2237 => "0000000000000000",
        2238 => "0000000000000000",
        2239 => "0000000000000000",
        2240 => "0000000000000000",
        2241 => "0000000000000000",
        2242 => "0000000000000000",
        2243 => "0000000000000000",
        2244 => "0000000000000000",
        2245 => "0000000000000000",
        2246 => "0000000000000000",
        2247 => "0000000000000000",
        2248 => "0000000000000000",
        2249 => "0000000000000000",
        2250 => "0000000000000000",
        2251 => "0000000000000000",
        2252 => "0000000000000000",
        2253 => "0000000000000000",
        2254 => "0000000000000000",
        2255 => "0000000000000000",
        2256 => "0000000000000000",
        2257 => "0000000000000000",
        2258 => "0000000000000000",
        2259 => "0000000000000000",
        2260 => "0000000000000000",
        2261 => "0000000000000000",
        2262 => "0000000000000000",
        2263 => "0000000000000000",
        2264 => "0000000000000000",
        2265 => "0000000000000000",
        2266 => "0000000000000000",
        2267 => "0000000000000000",
        2268 => "0000000000000000",
        2269 => "0000000000000000",
        2270 => "0000000000000000",
        2271 => "0000000000000000",
        2272 => "0000000000000000",
        2273 => "0000000000000000",
        2274 => "0000000000000000",
        2275 => "0000000000000000",
        2276 => "0000000000000000",
        2277 => "0000000000000000",
        2278 => "0000000000000000",
        2279 => "0000000000000000",
        2280 => "0000000000000000",
        2281 => "0000000000000000",
        2282 => "0000000000000000",
        2283 => "0000000000000000",
        2284 => "0000000000000000",
        2285 => "0000000000000000",
        2286 => "0000000000000000",
        2287 => "0000000000000000",
        2288 => "0000000000000000",
        2289 => "0000000000000000",
        2290 => "0000000000000000",
        2291 => "0000000000000000",
        2292 => "0000000000000000",
        2293 => "0000000000000000",
        2294 => "0000000000000000",
        2295 => "0000000000000000",
        2296 => "0000000000000000",
        2297 => "0000000000000000",
        2298 => "0000000000000000",
        2299 => "0000000000000000",
        2300 => "0000000000000000",
        2301 => "0000000000000000",
        2302 => "0000000000000000",
        2303 => "0000000000000000",
        2304 => "0000000000000000",
        2305 => "0000000000000000",
        2306 => "0000000000000000",
        2307 => "0000000000000000",
        2308 => "0000000000000000",
        2309 => "0000000000000000",
        2310 => "0000000000000000",
        2311 => "0000000000000000",
        2312 => "0000000000000000",
        2313 => "0000000000000000",
        2314 => "0000000000000000",
        2315 => "0000000000000000",
        2316 => "0000000000000000",
        2317 => "0000000000000000",
        2318 => "0000000000000000",
        2319 => "0000000000000000",
        2320 => "0000000000000000",
        2321 => "0000000000000000",
        2322 => "0000000000000000",
        2323 => "0000000000000000",
        2324 => "0000000000000000",
        2325 => "0000000000000000",
        2326 => "0000000000000000",
        2327 => "0000000000000000",
        2328 => "0000000000000000",
        2329 => "0000000000000000",
        2330 => "0000000000000000",
        2331 => "0000000000000000",
        2332 => "0000000000000000",
        2333 => "0000000000000000",
        2334 => "0000000000000000",
        2335 => "0000000000000000",
        2336 => "0000000000000000",
        2337 => "0000000000000000",
        2338 => "0000000000000000",
        2339 => "0000000000000000",
        2340 => "0000000000000000",
        2341 => "0000000000000000",
        2342 => "0000000000000000",
        2343 => "0000000000000000",
        2344 => "0000000000000000",
        2345 => "0000000000000000",
        2346 => "0000000000000000",
        2347 => "0000000000000000",
        2348 => "0000000000000000",
        2349 => "0000000000000000",
        2350 => "0000000000000000",
        2351 => "0000000000000000",
        2352 => "0000000000000000",
        2353 => "0000000000000000",
        2354 => "0000000000000000",
        2355 => "0000000000000000",
        2356 => "0000000000000000",
        2357 => "0000000000000000",
        2358 => "0000000000000000",
        2359 => "0000000000000000",
        2360 => "0000000000000000",
        2361 => "0000000000000000",
        2362 => "0000000000000000",
        2363 => "0000000000000000",
        2364 => "0000000000000000",
        2365 => "0000000000000000",
        2366 => "0000000000000000",
        2367 => "0000000000000000",
        2368 => "0000000000000000",
        2369 => "0000000000000000",
        2370 => "0000000000000000",
        2371 => "0000000000000000",
        2372 => "0000000000000000",
        2373 => "0000000000000000",
        2374 => "0000000000000000",
        2375 => "0000000000000000",
        2376 => "0000000000000000",
        2377 => "0000000000000000",
        2378 => "0000000000000000",
        2379 => "0000000000000000",
        2380 => "0000000000000000",
        2381 => "0000000000000000",
        2382 => "0000000000000000",
        2383 => "0000000000000000",
        2384 => "0000000000000000",
        2385 => "0000000000000000",
        2386 => "0000000000000000",
        2387 => "0000000000000000",
        2388 => "0000000000000000",
        2389 => "0000000000000000",
        2390 => "0000000000000000",
        2391 => "0000000000000000",
        2392 => "0000000000000000",
        2393 => "0000000000000000",
        2394 => "0000000000000000",
        2395 => "0000000000000000",
        2396 => "0000000000000000",
        2397 => "0000000000000000",
        2398 => "0000000000000000",
        2399 => "0000000000000000",
        2400 => "0000000000000000",
        2401 => "0000000000000000",
        2402 => "0000000000000000",
        2403 => "0000000000000000",
        2404 => "0000000000000000",
        2405 => "0000000000000000",
        2406 => "0000000000000000",
        2407 => "0000000000000000",
        2408 => "0000000000000000",
        2409 => "0000000000000000",
        2410 => "0000000000000000",
        2411 => "0000000000000000",
        2412 => "0000000000000000",
        2413 => "0000000000000000",
        2414 => "0000000000000000",
        2415 => "0000000000000000",
        2416 => "0000000000000000",
        2417 => "0000000000000000",
        2418 => "0000000000000000",
        2419 => "0000000000000000",
        2420 => "0000000000000000",
        2421 => "0000000000000000",
        2422 => "0000000000000000",
        2423 => "0000000000000000",
        2424 => "0000000000000000",
        2425 => "0000000000000000",
        2426 => "0000000000000000",
        2427 => "0000000000000000",
        2428 => "0000000000000000",
        2429 => "0000000000000000",
        2430 => "0000000000000000",
        2431 => "0000000000000000",
        2432 => "0000000000000000",
        2433 => "0000000000000000",
        2434 => "0000000000000000",
        2435 => "0000000000000000",
        2436 => "0000000000000000",
        2437 => "0000000000000000",
        2438 => "0000000000000000",
        2439 => "0000000000000000",
        2440 => "0000000000000000",
        2441 => "0000000000000000",
        2442 => "0000000000000000",
        2443 => "0000000000000000",
        2444 => "0000000000000000",
        2445 => "0000000000000000",
        2446 => "0000000000000000",
        2447 => "0000000000000000",
        2448 => "0000000000000000",
        2449 => "0000000000000000",
        2450 => "0000000000000000",
        2451 => "0000000000000000",
        2452 => "0000000000000000",
        2453 => "0000000000000000",
        2454 => "0000000000000000",
        2455 => "0000000000000000",
        2456 => "0000000000000000",
        2457 => "0000000000000000",
        2458 => "0000000000000000",
        2459 => "0000000000000000",
        2460 => "0000000000000000",
        2461 => "0000000000000000",
        2462 => "0000000000000000",
        2463 => "0000000000000000",
        2464 => "0000000000000000",
        2465 => "0000000000000000",
        2466 => "0000000000000000",
        2467 => "0000000000000000",
        2468 => "0000000000000000",
        2469 => "0000000000000000",
        2470 => "0000000000000000",
        2471 => "0000000000000000",
        2472 => "0000000000000000",
        2473 => "0000000000000000",
        2474 => "0000000000000000",
        2475 => "0000000000000000",
        2476 => "0000000000000000",
        2477 => "0000000000000000",
        2478 => "0000000000000000",
        2479 => "0000000000000000",
        2480 => "0000000000000000",
        2481 => "0000000000000000",
        2482 => "0000000000000000",
        2483 => "0000000000000000",
        2484 => "0000000000000000",
        2485 => "0000000000000000",
        2486 => "0000000000000000",
        2487 => "0000000000000000",
        2488 => "0000000000000000",
        2489 => "0000000000000000",
        2490 => "0000000000000000",
        2491 => "0000000000000000",
        2492 => "0000000000000000",
        2493 => "0000000000000000",
        2494 => "0000000000000000",
        2495 => "0000000000000000",
        2496 => "0000000000000000",
        2497 => "0000000000000000",
        2498 => "0000000000000000",
        2499 => "0000000000000000",
        2500 => "0000000000000000",
        2501 => "0000000000000000",
        2502 => "0000000000000000",
        2503 => "0000000000000000",
        2504 => "0000000000000000",
        2505 => "0000000000000000",
        2506 => "0000000000000000",
        2507 => "0000000000000000",
        2508 => "0000000000000000",
        2509 => "0000000000000000",
        2510 => "0000000000000000",
        2511 => "0000000000000000",
        2512 => "0000000000000000",
        2513 => "0000000000000000",
        2514 => "0000000000000000",
        2515 => "0000000000000000",
        2516 => "0000000000000000",
        2517 => "0000000000000000",
        2518 => "0000000000000000",
        2519 => "0000000000000000",
        2520 => "0000000000000000",
        2521 => "0000000000000000",
        2522 => "0000000000000000",
        2523 => "0000000000000000",
        2524 => "0000000000000000",
        2525 => "0000000000000000",
        2526 => "0000000000000000",
        2527 => "0000000000000000",
        2528 => "0000000000000000",
        2529 => "0000000000000000",
        2530 => "0000000000000000",
        2531 => "0000000000000000",
        2532 => "0000000000000000",
        2533 => "0000000000000000",
        2534 => "0000000000000000",
        2535 => "0000000000000000",
        2536 => "0000000000000000",
        2537 => "0000000000000000",
        2538 => "0000000000000000",
        2539 => "0000000000000000",
        2540 => "0000000000000000",
        2541 => "0000000000000000",
        2542 => "0000000000000000",
        2543 => "0000000000000000",
        2544 => "0000000000000000",
        2545 => "0000000000000000",
        2546 => "0000000000000000",
        2547 => "0000000000000000",
        2548 => "0000000000000000",
        2549 => "0000000000000000",
        2550 => "0000000000000000",
        2551 => "0000000000000000",
        2552 => "0000000000000000",
        2553 => "0000000000000000",
        2554 => "0000000000000000",
        2555 => "0000000000000000",
        2556 => "0000000000000000",
        2557 => "0000000000000000",
        2558 => "0000000000000000",
        2559 => "0000000000000000",
        2560 => "0000000000000000",
        2561 => "0010100000100000",
        2562 => "1111100000000000",
        others => (others => '0')
    );

    signal instruction_reg: std_logic_vector(15 downto 0); -- Register for instruction output
begin

    process(clk)
    begin
    -- write then read
        if rising_edge(clk) then
            if write_enable = '1' then
                memory(to_integer(unsigned(write_address))) <= write_data;
            end if;
        end if;
    end process;

    instruction_reg <= memory(to_integer(unsigned(pc))) when to_integer(unsigned(pc)) < 4096 else (others => '0');

    -- Output the instruction
    instruction <= instruction_reg;
end Behavioral;
